
///////////////////////////VIRTUAL INTERFACE
interface ram_if();
  logic clk;
  logic wr;
  logic [7:0] din;
  logic [7:0] dout;
  logic [3:0] addr;
endinterface
