interface intf(input bit clk);
  logic [2:0] Op_code;
  logic [31:0] A,B,Y;
endinterface